`ifndef TEST_BASE_SV
 `define TEST_BASE_SV

class test_base extends uvm_test;

   log_env env;
   log_config cfg;
   
   `uvm_component_utils(test_base)   
   
   function new(string name = "test_base", uvm_component parent = null);
      super.new(name,parent);
   endfunction : new

   function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      cfg = log_config::type_id::create("cfg");
      uvm_config_db#(log_config)::set(this,"env","log_config",cfg);
      env = log_env::type_id::create("env",this);
   endfunction : build_phase

   function void end_of_elaboration_phase(uvm_phase phase);
      super.end_of_elaboration_phase(phase);
      uvm_top.print_topology();
   endfunction: end_of_elaboration_phase

   function void init_vseq(virtual_seq vseq, virtual_seq1 vseq1, virtual_seq2 vseq2);
      vseq.sequencer_lite_if = env.agent.seqr;
      vseq1.sequencer_full_if = env.agent1.seqr1;
      vseq2.sequencer_lite1_if = env.agent.seqr;
   endfunction:init_vseq
  
   
endclass : test_base
`endif
